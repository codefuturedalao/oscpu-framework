`include "defines.v"
module encoder32_5(
        input [31 : 0] in,
        output [4 : 0] out

);
    assign out = ({5{in[0]}} & 5'b00000)
            |    ({5{in[1]}} & 5'b00001)
            |    ({5{in[2]}} & 5'b00010)
            |    ({5{in[3]}} & 5'b00011)
            |    ({5{in[4]}} & 5'b00100)
            |    ({5{in[5]}} & 5'b00101)
            |    ({5{in[6]}} & 5'b00110)
            |    ({5{in[7]}} & 5'b00111)
            |    ({5{in[8]}} & 5'b01000)
            |    ({5{in[9]}} & 5'b01001)
            |    ({5{in[10]}} & 5'b01010)
            |    ({5{in[11]}} & 5'b01011)
            |    ({5{in[12]}} & 5'b01100)
            |    ({5{in[13]}} & 5'b01101)
            |    ({5{in[14]}} & 5'b01110)
            |    ({5{in[15]}} & 5'b01111)
            |    ({5{in[16]}} & 5'b10000)
            |    ({5{in[17]}} & 5'b10001)
            |    ({5{in[18]}} & 5'b10010)
            |    ({5{in[19]}} & 5'b10011)
            |    ({5{in[20]}} & 5'b10100)
            |    ({5{in[21]}} & 5'b10101)
            |    ({5{in[22]}} & 5'b10110)
            |    ({5{in[23]}} & 5'b10111)
            |    ({5{in[24]}} & 5'b11000)
            |    ({5{in[25]}} & 5'b11001)
            |    ({5{in[26]}} & 5'b11010)
            |    ({5{in[27]}} & 5'b11011)
            |    ({5{in[28]}} & 5'b11100)
            |    ({5{in[29]}} & 5'b11101)
            |    ({5{in[30]}} & 5'b11110)
            |    ({5{in[31]}} & 5'b11111);

endmodule